`timescale 1ns/1ns
/*ģ��˵��
����һ��ʱ��ģ�飬���ʱ���룬���밴��
key4�������ã��ͼ�ʱ��״̬�л�
������״̬�£�key1,2,3�ֱ����ʱ���룬��һ�£���һ��
*/
module clock (
    //global clock
    input        clk,
    input        rst_n,

    //user interface
    input  [3:0] key,

    output [7:0] hour,
    output [7:0] minu,
    output [7:0] seco
);

wire rst;

reg [25:0]cnt0;
wire add_cnt0;
wire end_cnt0;
reg [5:0]cnt1;
wire add_cnt1;
wire end_cnt1;
reg [5:0]cnt2;
wire add_cnt2;
wire end_cnt2;
reg [5:0]cnt3;
wire add_cnt3;
wire end_cnt3;

reg [1:0] state_c, state_n;
wire set_to_tim_start ;
wire tim_to_set_start ;


localparam  set = 1;
localparam  tim = 2;

rst rst_u(
    //global clock
    . clk(clk),
    . rst_n(rst_n),

    //user interface
    . rst(rst)
);

assign seco = {(cnt1/10)%10,cnt1%10};
assign hour = 0;
assign minu = 0;
always @(posedge clk or negedge rst) begin
    if (!rst_n)
        state_c <= set ;
    else
        state_c <= state_n;
end

always @(*) begin
    case(state_c)
        set :begin
            if(set_to_tim_start)
                state_n = tim ;
            else
                state_n = state_c ;
        end
        tim :begin
            if(tim_to_set_start)
                state_n = set ;
            else
                state_n = state_c ;
        end
        default : state_n = set ;
    endcase
end

assign set_to_tim_start = state_c==set && (key[3]);
assign tim_to_set_start = state_c==tim && (key[3]);



//������0 seco
    always @(posedge clk or negedge rst)begin
        if(!rst_n)begin
            cnt0 <= 0;
          end
        else if(add_cnt0)begin
          if(end_cnt0)
             cnt0 <= 0;
          else 
             cnt0 <= cnt0 + 1;
          end      
    end

assign add_cnt0 = state_c == tim;
assign end_cnt0 = add_cnt0 && cnt0 == 50_0-1;//50_000_000-1

//������1 minu
    always @(posedge clk or negedge rst)begin
        if(!rst_n)begin
            cnt1 <= 0;
          end
        else if(add_cnt1)begin
          if(end_cnt1)
             cnt1 <= 0; 
          else
             cnt1 <= cnt1 + 1; 
        end
    end

assign add_cnt1 = end_cnt0 || key[2] == 1;
assign end_cnt1 = add_cnt1 && cnt1 == 60-1;

//������2 hour
    always @(posedge clk or negedge rst)begin
        if(!rst_n)begin
            cnt2 <= 0;
          end
        else if(add_cnt2)begin
          if(end_cnt2)
             cnt2 <= 0;
          else
             cnt2 <= cnt2 + 1;     
        end
    end

assign add_cnt2 = end_cnt1 || key[1] == 1;
assign end_cnt2 = add_cnt2 && cnt2 == 60-1;

//������3 day
    always @(posedge clk or negedge rst)begin
        if(!rst_n)begin
            cnt3 <= 0;
          end
        else if(add_cnt3)begin
          if(end_cnt3)
             cnt3 <= 0;
          else
             cnt3 <= cnt3 + 1;     
        end
    end

assign add_cnt3 = end_cnt2 || key[0] == 1;
assign end_cnt3 = add_cnt3 && cnt3 == 24-1;
    
endmodule